`timescale 1ns / 1ps
`include "macro.vh"

// `define LEN1 (16)
// `define LEN2 (16)
// `define MAX_LEN1 (16)
// `define MAX_LEN2 (16)

`define MAX_LEN1 (1024)
`define MAX_LEN2 (1536)
`define PIPELINE_LENGTH (48)


import datatypesPkg::*;

module tb_med_solver_with_ram(output logic finished, output logic grid_finished,
            output logic [$clog2(`MAX_LEN1):0] maxRowId,
            output logic [$clog2(`MAX_LEN2):0] maxColId,
            output logic [0:`MAX_LEN1-1] [15:0] score_grid [0:192-1],
            output direction grid [0:`PIPELINE_LENGTH-1] [0:(`MAX_LEN1*`MAX_LEN2/`PIPELINE_LENGTH)-1],
            output direction aligned_sequence [0:`MAX_LEN1+`MAX_LEN2-1]
);

    logic clk;      // clock signal we are going to generate
    logic rst;      // the reset input used to initialise the system
    logic solver_enable;

    // dna_base seq1 [`MAX_LEN1-1:0] = '{A,T,C,A,G,T,A,T,C,A,G,T,T,G,G, A};
    // dna_base seq2 [`MAX_LEN2-1:0] = '{G,G,C,A,G,G,C,A,G,G,C,T,T,G,T, A};

    // dna_base seq1 [0:`MAX_LEN1-1] = '{A ,G,T,T,G,A,C,T,A,T,G,A,C,T,A,C,G,G,T,T,G,A,C,T,A,T,G,A,C,T,A,C,G,G,T,T,G,A,C,T,A,T,G,A,C,T,A,C,G,G,T,T,G,A,C,T,A,T,G,A,C,T,A,C, A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A,A};
    // dna_base seq2 [0:`MAX_LEN2-1] = '{A ,A,G,G,C,G,A,C,G,G,C,T,G,T,T,C,G,G,A,C,G,G,A,C,T,G,T,T,C,G,G,A,C,G,G,A,C,G,G,C,T,G,T,G,T,T,C,G,G,A,C,G,G,T,T,C,G,G,A,C,G,G,G,C};

    `seq_base seq1 [0:`MAX_LEN1-1]; // = '{A, A,G,G,G,G,C,G,T,T,G,T,A,G,A,T,C,T,C,T,C,A,G,C,C,C,T,G,A,T,G,T,A,G,G,G,G,G,C,C,G,C,A,G,C,A,A,C,G,C,T,C,T,G,T,T,T,G,T,G,A,C,G,T,A,T,G,T,T,G,T,T,G,T,C,T,C,T,A,T,C,C,A,A,C,C,C,C,G,G,C,C,C,T,A,T,A,A,A,T,T,T,T,T,G,A,G,A,T,G,T,C,C,G,A,C,G,A,C,C,G,G,T,C,A,G,A,A,A,T,C,C,T,G,G,T,T,C,A,G,C,G,C,A,A,A,A,G,G,T,C,A,C,T,T,A,A,G,A,T,C,A,A,A,G,A,A,G,G,G,G,C,A,C,C,A,T,C,C,G,A,G,T,T,T,C,C,C,T,T,C,T,G,A,A,G,T,A,G,T,T,C,T,T,C,C,A,G,A,T,C,T,T,C,T,T,G,C,T,C,C,G,A,C,A,T,A,C,A,G,T,C,G,A,A,G,G,G,A,T,A,A,T,A,C,C,A,T,C,A,A,C,T,A,G,C,G,T,C,A,A,C,T,C,A,A,C,T,C,A,C,T,G,G,T,A,G,T,T,C,C,T,G,C,T,G,A,G,A,A,T,A,C,T,T,T,A,T,A,T,G,T,G,A,A,A,T,G,G,C,A,T,G,C,C,A,T,A,G,T,A,C,T,G,C,A,C,C,A,A,G,C,G,C,T,G,A,A,T,T,A,G,T,A,T,C,G,G,A,T,G,G,T,A,T,T,C,A,G,C,A,T,G,C,C,T,A,A,A,G,G,C,A,T,G,G,G,T,T,A,C,C,T,C,G,C,C,C,G,G,T,T,A,C,C,T,A,C,G,C,A,T,T,A,G,A,C,T,G,G,T,C,A,T,A,G,A,C,C,C,C,G,T,A,T,T,A,T,C,T,T,T,T,C,T,C,T,G,G,G,C,C,A,C,G,C,A,G,G,C,T,G,T,T,C,A,C,C,G,C,T,G,A,G,C,G,G,T,C,G,A,C,A,C,C,G,A,T,G,C,T,G,G,A,G,G,G,T,T,G,C,G,A,G,C,A,C,G,T,A,G,C,A,G,G,C,A,T,C,A,T,C,T,G,G,A,C,A,G,T,G,G,G,T,A,A,G,A,T,T,A,C,G,G,C,T,T,A,A,T,T,G,T,A,T,C,G,C,G,T,C,G,G,A,A,C,G,A,A,C,A,A,G,G,T,G,C,A,G,C,A,T,A,T,C,C,G,T,A,A,T,T,T,T,C,T,C,C,A,A,A,T,C,G,C,A,C,C,A,T,T,G,G,A,A,C,A,G,C,T,A,A,A,G,T,G,A,G,A,G,A,A,C,C,G,T,A,G,G,T,A,T,C,C,C,T,C,A,C,G,G,A,C,C,G,C,C,A,C,C,A,A,A,T,C,A,A,A,A,C,C,T,T,A,A,A,C,G,T,A,T,G,G,C,A,T,T,A,G,G,C,T,A,A,C,C,A,C,A,C,T,T,A,G,T,C,A,T,G,G,C,C,G,C,G,T,T,C,C,T,G,G,A,C,G,A,G,G,G,A,C,G,G,A,A,A,T,T,A,A,G,G,G,C,C,G,T,G,G,A,G,G,G,A,C,C,C,T,G,G,C,G,A,C,A,G,G,T,C,T,A,A,C,G,G,G,T,G,T,T,C,C,T,A,T,A,T,C,C,A,A,C,C,T,C,T,A,G,C,A,T,C,C,C,T,A,C,A,C,G,T,A,G,A,C,C,T,C,A,A,T,G,A,G,C,G,G,T,G,C,G,C,A,A,G,A,T,T,T,G,C,C,C,T,T,A,G,A,T,G,T,G,C,G,C,T,C,A,T,G,C,T,T,T,G,T,C,T,T,T,A,G,A,C,C,C,C,G,A,A,C,T,C,T,G,C,A,G,G,C,T,C,C,A,C,A,T,C,T,G,T,T,T,C,A,C,G,A,T,A,A,A,T,C,C,C,A,G,C,G,T,C,T,A,T,G,A,T,G,T,G,G,T,A,G,C,G,T,C,C,C,G,T,C,A,T,C,T,A,T,T,A,C,G,G,T,A,A,T,G,G,C,C,G,T,T,A,T,G,A,A,T,G,T,C,T,T,A,T,G,C,T,G,C,C,G,A,G,C,T,T,C,T,G,G,A,C,G,A,G,T,C,T,A,G,T,C,T,C,C,T,A,T,A,G,T,A,T,G,G,G,A,C,G,G,G,C,T,C,T,G,A,C,T};
    `seq_base seq2 [0:`MAX_LEN2-1]; // = '{A, G,A,C,C,T,T,A,C,G,T,C,A,C,C,T,T,T,G,C,A,T,C,T,C,G,A,C,G,A,A,T,T,T,C,G,A,T,C,G,A,C,C,A,T,G,G,A,T,A,T,T,C,T,T,G,C,T,G,C,G,T,C,T,T,C,A,G,A,G,T,T,G,C,C,A,T,G,G,A,C,G,G,G,G,A,A,C,G,A,G,T,G,G,A,T,A,C,A,C,C,T,C,C,C,G,A,C,T,T,T,A,A,A,C,A,G,A,A,A,T,C,G,T,C,G,C,A,T,A,C,T,C,T,G,C,C,T,A,T,C,G,C,A,C,T,C,T,T,G,A,C,T,A,C,A,T,G,G,T,G,G,G,G,A,C,T,C,C,T,T,A,T,C,A,G,C,T,C,G,A,C,T,T,G,G,G,G,C,C,C,A,A,G,G,T,A,C,A,A,G,T,A,G,G,T,T,G,A,A,A,C,G,G,C,C,C,G,G,C,G,T,T,G,T,T,G,G,C,G,T,C,A,C,T,C,T,T,A,G,C,A,C,A,C,T,G,A,C,G,C,T,C,C,T,A,G,C,T,G,A,G,A,C,C,T,T,G,A,A,C,A,T,G,C,A,G,G,A,C,G,T,C,C,C,T,G,T,G,C,C,A,A,T,T,C,G,C,T,A,T,G,G,G,C,C,T,T,C,A,A,G,G,A,T,T,T,C,A,T,A,G,C,A,T,T,A,C,C,G,T,C,T,C,A,C,G,G,C,C,A,C,G,C,A,G,G,G,C,G,C,G,A,T,G,A,A,C,C,C,G,G,T,T,A,G,T,T,G,A,T,T,T,T,G,T,G,A,T,T,T,A,T,T,T,C,G,T,G,T,G,G,T,C,A,T,A,C,G,C,G,G,A,T,T,C,T,T,A,C,T,A,A,G,T,C,T,C,T,A,C,G,G,A,A,G,A,A,C,C,C,T,C,G,A,T,A,G,G,A,G,T,C,C,G,A,C,A,A,T,G,G,A,G,A,A,T,A,A,C,T,A,A,A,G,A,A,G,C,G,C,T,T,C,G,A,C,C,C,C,A,A,G,C,G,A,C,A,G,C,G,A,A,T,C,G,G,G,A,T,T,T,G,C,G,A,G,A,A,C,T,C,A,C,A,G,G,A,T,C,C,A,T,C,A,A,G,T,C,C,T,A,C,C,G,T,C,G,C,T,G,A,G,C,A,G,G,T,C,C,T,G,G,G,A,C,A,G,T,A,G,T,T,C,C,A,G,T,T,A,T,T,C,C,T,A,A,T,A,G,A,C,T,C,A,G,C,T,C,C,A,G,C,A,G,G,A,G,C,G,A,C,T,A,A,A,A,G,G,T,C,A,A,A,G,G,G,A,C,C,T,C,T,T,G,G,G,G,T,T,G,A,G,C,G,A,C,C,T,G,T,G,T,T,T,T,A,A,C,G,C,C,A,G,G,C,C,C,T,A,A,C,C,C,C,G,C,C,T,G,G,A,G,G,G,C,C,C,G,C,A,A,G,T,G,G,T,C,A,G,C,T,G,T,T,C,T,A,G,T,A,C,A,G,T,T,A,C,T,G,A,T,C,A,G,A,A,T,C,A,C,T,G,T,C,C,G,C,C,T,A,C,C,C,G,T,T,C,A,T,C,C,A,A,C,G,T,G,G,T,T,T,G,A,C,G,A,T,T,C,C,C,G,A,G,G,G,T,A,A,T,A,T,A,G,G,C,C,G,G,C,A,C,T,A,T,T,C,G,C,G,G,C,G,T,T,A,G,T,T,G,T,T,C,T,T,C,C,T,G,C,C,G,G,A,C,A,C,C,T,A,T,C,C,T,C,G,A,C,T,C,G,G,C,G,C,G,G,G,G,A,G,C,C,A,G,A,A,C,G,C,G,A,T,G,T,G,T,G,A,A,C,T,T,C,G,G,T,C,C,G,G,C,A,A,A,A,A,A,A,C,C,A,T,A,T,C,G,T,G,G,T,A,C,C,G,C,T,A,G,T,A,A,T,C,A,C,T,T,C,T,A,G,T,T,T,C,T,G,T,G,A,A,G,T,C,G,G,A,C,T,C,C,G,A,T,C,C,G,A,A,C,C,A,A,G,A,G,T,A,C,G,G,A,G,A,A,T,T,C,G,A,A,G,C,G,C,T,G,C,C,G,A,T,G,C,A,C,T,C,G,C,C,A,G,A,G,G,T,A,G,C,C,G,C,A,C,T,A,A,T,A,T,C,C,G,G,T,G,A,A,C,A,G,G,T,A,G,T,G,C,G,A,G};

    logic [11:0] len1;
    logic [12:0] len2;

    logic rdreq;
    logic wrreq;
    logic sclr;

    logic empty;
    logic full;

    logic [15:0] in16;
    logic [15:0] out16;

    logic [1:0] in2;
    logic [1:0] out2;
    logic [14:0] wraddress;
    logic [14:0] rdaddress;
    logic wren;

                    // instantiate design under test
    fifo_16b_1024w last_col (.aclr(rst), .clock(clk), .sclr(sclr),
        .data(in16), .rdreq(rdreq),
        .q(out16), .wrreq(wrreq),
        .empty(empty), .full(full)
    );

    pe_bram pe_cell_bram (
        .data(in2),
        .rdaddress(rdaddress),
        .rdclock(clk),
        .rd_aclr(rst),
        .wraddress(wraddress),
        .wrclock(clk),
        .wren(wren),
        .q(out2)
    );


    med_solver_with_ram #(.max_len1(`MAX_LEN1), .max_len2(`MAX_LEN2), .pipeline_length(`PIPELINE_LENGTH)) ms
    (.clk(clk), .rst(rst), .solver_enable(solver_enable), .len1(len1), .len2(len2), .seq1(seq1), .seq2(seq2),
    .finished(finished), .grid_finished(grid_finished), .maxRowId(maxRowId), .maxColId(maxColId),
    // .grid(grid), .score_grid(score_grid),
    .aligned_sequence(aligned_sequence));


    initial          // sequence of events to simulate
        begin
            clk = 0;     // at time=0 set clock to zero and reset to active (1)
            rst = 1;
            solver_enable = 0;

            sclr = 1'b0;
            rdreq = 1'b0;
            wrreq = 1'b0;
            in16 = 16'hFF00;

            wren = 1'b0;
            in2 = 2'b11;
            rdaddress = 15'd2;
            wraddress = 15'd2;

            seq1 = '{nA, nA,nG,nG,nG,nG,nC,nG,nT,nT,nG,nT,nA,nG,nA,nT,nC,nT,nC,nT,nC,nA,nG,nC,nC,nC,nT,nG,nA,nT,nG,nT,nA,nG,nG,nG,nG,nG,nC,nC,nG,nC,nA,nG,nC,nA,nA,nC,nG,nC,nT,nC,nT,nG,nT,nT,nT,nG,nT,nG,nA,nC,nG,nT,nA,nT,nG,nT,nT,nG,nT,nT,nG,nT,nC,nT,nC,nT,nA,nT,nC,nC,nA,nA,nC,nC,nC,nC,nG,nG,nC,nC,nC,nT,nA,nT,nA,nA,nA,nT,nT,nT,nT,nT,nG,nA,nG,nA,nT,nG,nT,nC,nC,nG,nA,nC,nG,nA,nC,nC,nG,nG,nT,nC,nA,nG,nA,nA,nA,nT,nC,nC,nT,nG,nG,nT,nT,nC,nA,nG,nC,nG,nC,nA,nA,nA,nA,nG,nG,nT,nC,nA,nC,nT,nT,nA,nA,nG,nA,nT,nC,nA,nA,nA,nG,nA,nA,nG,nG,nG,nG,nC,nA,nC,nC,nA,nT,nC,nC,nG,nA,nG,nT,nT,nT,nC,nC,nC,nT,nT,nC,nT,nG,nA,nA,nG,nT,nA,nG,nT,nT,nC,nT,nT,nC,nC,nA,nG,nA,nT,nC,nT,nT,nC,nT,nT,nG,nC,nT,nC,nC,nG,nA,nC,nA,nT,nA,nC,nA,nG,nT,nC,nG,nA,nA,nG,nG,nG,nA,nT,nA,nA,nT,nA,nC,nC,nA,nT,nC,nA,nA,nC,nT,nA,nG,nC,nG,nT,nC,nA,nA,nC,nT,nC,nA,nA,nC,nT,nC,nA,nC,nT,nG,nG,nT,nA,nG,nT,nT,nC,nC,nT,nG,nC,nT,nG,nA,nG,nA,nA,nT,nA,nC,nT,nT,nT,nA,nT,nA,nT,nG,nT,nG,nA,nA,nA,nT,nG,nG,nC,nA,nT,nG,nC,nC,nA,nT,nA,nG,nT,nA,nC,nT,nG,nC,nA,nC,nC,nA,nA,nG,nC,nG,nC,nT,nG,nA,nA,nT,nT,nA,nG,nT,nA,nT,nC,nG,nG,nA,nT,nG,nG,nT,nA,nT,nT,nC,nA,nG,nC,nA,nT,nG,nC,nC,nT,nA,nA,nA,nG,nG,nC,nA,nT,nG,nG,nG,nT,nT,nA,nC,nC,nT,nC,nG,nC,nC,nC,nG,nG,nT,nT,nA,nC,nC,nT,nA,nC,nG,nC,nA,nT,nT,nA,nG,nA,nC,nT,nG,nG,nT,nC,nA,nT,nA,nG,nA,nC,nC,nC,nC,nG,nT,nA,nT,nT,nA,nT,nC,nT,nT,nT,nT,nC,nT,nC,nT,nG,nG,nG,nC,nC,nA,nC,nG,nC,nA,nG,nG,nC,nT,nG,nT,nT,nC,nA,nC,nC,nG,nC,nT,nG,nA,nG,nC,nG,nG,nT,nC,nG,nA,nC,nA,nC,nC,nG,nA,nT,nG,nC,nT,nG,nG,nA,nG,nG,nG,nT,nT,nG,nC,nG,nA,nG,nC,nA,nC,nG,nT,nA,nG,nC,nA,nG,nG,nC,nA,nT,nC,nA,nT,nC,nT,nG,nG,nA,nC,nA,nG,nT,nG,nG,nG,nT,nA,nA,nG,nA,nT,nT,nA,nC,nG,nG,nC,nT,nT,nA,nA,nT,nT,nG,nT,nA,nT,nC,nG,nC,nG,nT,nC,nG,nG,nA,nA,nC,nG,nA,nA,nC,nA,nA,nG,nG,nT,nG,nC,nA,nG,nC,nA,nT,nA,nT,nC,nC,nG,nT,nA,nA,nT,nT,nT,nT,nC,nT,nC,nC,nA,nA,nA,nT,nC,nG,nC,nA,nC,nC,nA,nT,nT,nG,nG,nA,nA,nC,nA,nG,nC,nT,nA,nA,nA,nG,nT,nG,nA,nG,nA,nG,nA,nA,nC,nC,nG,nT,nA,nG,nG,nT,nA,nT,nC,nC,nC,nT,nC,nA,nC,nG,nG,nA,nC,nC,nG,nC,nC,nA,nC,nC,nA,nA,nA,nT,nC,nA,nA,nA,nA,nC,nC,nT,nT,nA,nA,nA,nC,nG,nT,nA,nT,nG,nG,nC,nA,nT,nT,nA,nG,nG,nC,nT,nA,nA,nC,nC,nA,nC,nA,nC,nT,nT,nA,nG,nT,nC,nA,nT,nG,nG,nC,nC,nG,nC,nG,nT,nT,nC,nC,nT,nG,nG,nA,nC,nG,nA,nG,nG,nG,nA,nC,nG,nG,nA,nA,nA,nT,nT,nA,nA,nG,nG,nG,nC,nC,nG,nT,nG,nG,nA,nG,nG,nG,nA,nC,nC,nC,nT,nG,nG,nC,nG,nA,nC,nA,nG,nG,nT,nC,nT,nA,nA,nC,nG,nG,nG,nT,nG,nT,nT,nC,nC,nT,nA,nT,nA,nT,nC,nC,nA,nA,nC,nC,nT,nC,nT,nA,nG,nC,nA,nT,nC,nC,nC,nT,nA,nC,nA,nC,nG,nT,nA,nG,nA,nC,nC,nT,nC,nA,nA,nT,nG,nA,nG,nC,nG,nG,nT,nG,nC,nG,nC,nA,nA,nG,nA,nT,nT,nT,nG,nC,nC,nC,nT,nT,nA,nG,nA,nT,nG,nT,nG,nC,nG,nC,nT,nC,nA,nT,nG,nC,nT,nT,nT,nG,nT,nC,nT,nT,nT,nA,nG,nA,nC,nC,nC,nC,nG,nA,nA,nC,nT,nC,nT,nG,nC,nA,nG,nG,nC,nT,nC,nC,nA,nC,nA,nT,nC,nT,nG,nT,nT,nT,nC,nA,nC,nG,nA,nT,nA,nA,nA,nT,nC,nC,nC,nA,nG,nC,nG,nT,nC,nT,nA,nT,nG,nA,nT,nG,nT,nG,nG,nT,nA,nG,nC,nG,nT,nC,nC,nC,nG,nT,nC,nA,nT,nC,nT,nA,nT,nT,nA,nC,nG,nG,nT,nA,nA,nT,nG,nG,nC,nC,nG,nT,nT,nA,nT,nG,nA,nA,nT,nG,nT,nC,nT,nT,nA,nT,nG,nC,nT,nG,nC,nC,nG,nA,nG,nC,nT,nT,nC,nT,nG,nG,nA,nC,nG,nA,nG,nT,nC,nT,nA,nG,nT,nC,nT,nC,nC,nT,nA,nT,nA,nG,nT,nA,nT,nG,nG,nG,nA,nC,nG,nG,nG,nC,nT,nC,nT,nG,nA,nC,nT};
            seq2 = '{nA, nG,nA,nC,nC,nT,nT,nA,nC,nG,nT,nC,nA,nC,nC,nT,nT,nT,nG,nC,nA,nT,nC,nT,nC,nG,nA,nC,nG,nA,nA,nT,nT,nT,nC,nG,nA,nT,nC,nG,nA,nC,nC,nA,nT,nG,nG,nA,nT,nA,nT,nT,nC,nT,nT,nG,nC,nT,nG,nC,nG,nT,nC,nT,nT,nC,nA,nG,nA,nG,nT,nT,nG,nC,nC,nA,nT,nG,nG,nA,nC,nG,nG,nG,nG,nA,nA,nC,nG,nA,nG,nT,nG,nG,nA,nT,nA,nC,nA,nC,nC,nT,nC,nC,nC,nG,nA,nC,nT,nT,nT,nA,nA,nA,nC,nA,nG,nA,nA,nA,nT,nC,nG,nT,nC,nG,nC,nA,nT,nA,nC,nT,nC,nT,nG,nC,nC,nT,nA,nT,nC,nG,nC,nA,nC,nT,nC,nT,nT,nG,nA,nC,nT,nA,nC,nA,nT,nG,nG,nT,nG,nG,nG,nG,nA,nC,nT,nC,nC,nT,nT,nA,nT,nC,nA,nG,nC,nT,nC,nG,nA,nC,nT,nT,nG,nG,nG,nG,nC,nC,nC,nA,nA,nG,nG,nT,nA,nC,nA,nA,nG,nT,nA,nG,nG,nT,nT,nG,nA,nA,nA,nC,nG,nG,nC,nC,nC,nG,nG,nC,nG,nT,nT,nG,nT,nT,nG,nG,nC,nG,nT,nC,nA,nC,nT,nC,nT,nT,nA,nG,nC,nA,nC,nA,nC,nT,nG,nA,nC,nG,nC,nT,nC,nC,nT,nA,nG,nC,nT,nG,nA,nG,nA,nC,nC,nT,nT,nG,nA,nA,nC,nA,nT,nG,nC,nA,nG,nG,nA,nC,nG,nT,nC,nC,nC,nT,nG,nT,nG,nC,nC,nA,nA,nT,nT,nC,nG,nC,nT,nA,nT,nG,nG,nG,nC,nC,nT,nT,nC,nA,nA,nG,nG,nA,nT,nT,nT,nC,nA,nT,nA,nG,nC,nA,nT,nT,nA,nC,nC,nG,nT,nC,nT,nC,nA,nC,nG,nG,nC,nC,nA,nC,nG,nC,nA,nG,nG,nG,nC,nG,nC,nG,nA,nT,nG,nA,nA,nC,nC,nC,nG,nG,nT,nT,nA,nG,nT,nT,nG,nA,nT,nT,nT,nT,nG,nT,nG,nA,nT,nT,nT,nA,nT,nT,nT,nC,nG,nT,nG,nT,nG,nG,nT,nC,nA,nT,nA,nC,nG,nC,nG,nG,nA,nT,nT,nC,nT,nT,nA,nC,nT,nA,nA,nG,nT,nC,nT,nC,nT,nA,nC,nG,nG,nA,nA,nG,nA,nA,nC,nC,nC,nT,nC,nG,nA,nT,nA,nG,nG,nA,nG,nT,nC,nC,nG,nA,nC,nA,nA,nT,nG,nG,nA,nG,nA,nA,nT,nA,nA,nC,nT,nA,nA,nA,nG,nA,nA,nG,nC,nG,nC,nT,nT,nC,nG,nA,nC,nC,nC,nC,nA,nA,nG,nC,nG,nA,nC,nA,nG,nC,nG,nA,nA,nT,nC,nG,nG,nG,nA,nT,nT,nT,nG,nC,nG,nA,nG,nA,nA,nC,nT,nC,nA,nC,nA,nG,nG,nA,nT,nC,nC,nA,nT,nC,nA,nA,nG,nT,nC,nC,nT,nA,nC,nC,nG,nT,nC,nG,nC,nT,nG,nA,nG,nC,nA,nG,nG,nT,nC,nC,nT,nG,nG,nG,nA,nC,nA,nG,nT,nA,nG,nT,nT,nC,nC,nA,nG,nT,nT,nA,nT,nT,nC,nC,nT,nA,nA,nT,nA,nG,nA,nC,nT,nC,nA,nG,nC,nT,nC,nC,nA,nG,nC,nA,nG,nG,nA,nG,nC,nG,nA,nC,nT,nA,nA,nA,nA,nG,nG,nT,nC,nA,nA,nA,nG,nG,nG,nA,nC,nC,nT,nC,nT,nT,nG,nG,nG,nG,nT,nT,nG,nA,nG,nC,nG,nA,nC,nC,nA,nC,nA,nG,nG,nA,nT,nC,nC,nA,nT,nC,nA,nA,nG,nT,nC,nC,nT,nA,nC,nC,nG,nT,nC,nG,nC,nT,nG,nA,nG,nC,nA,nG,nG,nT,nC,nC,nT,nG,nG,nG,nA,nC,nA,nG,nT,nA,nG,nT,nT,nC,nC,nA,nG,nT,nT,nA,nT,nT,nC,nC,nT,nA,nA,nT,nA,nG,nA,nC,nT,nC,nA,nG,nC,nT,nC,nC,nA,nG,nC,nA,nG,nG,nA,nG,nC,nG,nA,nC,nT,nA,nA,nA,nA,nG,nG,nT,nC,nA,nA,nA,nG,nG,nG,nA,nC,nC,nT,nC,nT,nT,nG,nG,nG,nG,nT,nT,nG,nA,nG,nC,nG,nA,nC,nC,nT,nG,nT,nG,nT,nT,nT,nT,nA,nA,nC,nG,nC,nC,nA,nG,nG,nC,nC,nC,nT,nA,nA,nC,nC,nC,nC,nG,nC,nC,nT,nG,nG,nA,nG,nG,nG,nC,nC,nC,nG,nC,nA,nA,nG,nT,nG,nG,nT,nC,nA,nG,nC,nT,nG,nT,nT,nC,nT,nA,nG,nT,nA,nC,nA,nG,nT,nT,nA,nC,nT,nG,nA,nT,nC,nA,nG,nA,nA,nT,nC,nA,nC,nT,nG,nT,nC,nC,nG,nC,nC,nT,nA,nC,nC,nC,nG,nT,nT,nC,nA,nT,nC,nC,nA,nA,nC,nG,nT,nG,nG,nT,nT,nT,nG,nA,nC,nG,nA,nT,nT,nC,nC,nC,nG,nA,nG,nG,nG,nT,nA,nA,nT,nA,nT,nA,nG,nG,nC,nC,nG,nG,nC,nA,nC,nT,nA,nT,nT,nC,nG,nC,nG,nG,nC,nG,nT,nT,nA,nG,nT,nT,nG,nT,nT,nC,nT,nT,nC,nC,nT,nG,nC,nC,nG,nG,nA,nC,nA,nC,nC,nT,nA,nT,nC,nC,nT,nC,nG,nA,nC,nT,nC,nG,nG,nC,nG,nC,nG,nG,nG,nG,nA,nG,nC,nC,nA,nG,nA,nA,nC,nG,nC,nG,nA,nT,nG,nT,nG,nT,nG,nA,nA,nC,nT,nT,nC,nG,nG,nT,nC,nC,nG,nG,nC,nA,nA,nA,nA,nA,nA,nA,nC,nC,nA,nT,nA,nT,nC,nG,nT,nG,nG,nT,nA,nC,nC,nG,nC,nT,nA,nG,nT,nA,nA,nT,nC,nA,nC,nT,nT,nC,nT,nA,nG,nT,nT,nT,nC,nT,nG,nT,nG,nA,nA,nG,nT,nC,nG,nG,nA,nC,nT,nC,nC,nG,nA,nT,nC,nC,nG,nA,nA,nC,nC,nA,nA,nG,nA,nG,nT,nA,nC,nG,nG,nA,nG,nA,nA,nT,nT,nC,nG,nA,nA,nG,nC,nG,nC,nT,nG,nC,nC,nG,nA,nT,nG,nC,nA,nC,nT,nC,nG,nC,nC,nA,nG,nA,nG,nG,nT,nA,nG,nC,nC,nG,nC,nA,nC,nT,nA,nA,nT,nA,nT,nC,nC,nG,nG,nT,nG,nA,nA,nC,nA,nG,nG,nT,nA,nG,nT,nG,nC,nG,nA,nG,nT,nG,nT,nG,nT,nT,nT,nT,nA,nA,nC,nG,nC,nC,nA,nG,nG,nC,nC,nC,nT,nA,nA,nC,nC,nC,nC,nG,nC,nC,nT,nG,nG,nA,nG,nG,nG,nC,nC,nC,nG,nC,nA,nA,nG,nT,nG,nG,nT,nC,nA,nG,nC,nT,nG,nT,nT,nC,nT,nA,nG,nT,nA,nC,nA,nG,nT,nT,nA,nC,nT,nG,nA,nT,nC,nA,nG,nA,nA,nT,nC,nA,nC,nT,nG,nT,nC,nC,nG,nC,nC,nT,nA,nC,nC,nC,nG,nT,nT,nC,nA,nT,nC,nC,nA,nA,nC,nG,nT,nG,nG,nT,nT,nT,nG,nA,nC,nG,nA,nT,nT,nC,nC,nC,nG,nA,nG,nG,nG,nT,nA,nA,nT,nA,nT,nA,nG,nG,nC,nC,nG,nG,nC,nA,nC,nT,nA,nT,nT,nC,nG,nC,nG,nG,nC,nG,nT,nT,nA,nG,nT,nT,nG,nT,nT,nC,nT,nT,nC,nC,nT,nG,nC,nC,nG,nG,nA,nC,nA,nC,nC,nT,nA,nT,nC,nC,nT,nC,nG,nA,nC,nT,nC,nG,nG,nC,nG,nC,nG,nG,nG,nG,nA,nG,nC,nC,nA,nG,nA,nA,nC,nG,nC,nG,nA,nT,nG,nT,nG,nT,nG,nA,nA,nC,nT,nT,nC,nG,nG,nT,nC,nC,nG,nG,nC,nA,nA,nA,nA,nA,nA,nA,nC,nC,nA,nT,nA,nT,nC,nG,nT,nG,nG,nT,nA,nC,nC,nG,nC,nT,nA,nG,nT,nA,nA,nT,nC,nA,nC,nT,nT,nC,nT,nA,nG,nT,nT,nT,nC,nT,nG,nT,nG,nA,nA,nG,nT,nC,nG,nG,nA,nC,nT,nC,nC,nG,nA,nT,nC,nC,nG,nA,nA,nC,nC,nA,nA,nG,nA,nG,nT,nA,nC,nG,nG,nA,nG,nA,nA,nT,nT,nC,nG,nA,nA,nG,nC,nG,nC,nT,nG,nC,nC,nG,nA,nT,nG,nC,nA,nC,nT,nC,nG,nC,nC,nA,nG,nA,nG,nG,nT,nA,nG,nC,nC,nG,nC,nA,nC,nT,nA,nA,nT,nA,nT,nC,nC,nG,nG,nT,nG,nA,nA,nC,nA,nG,nG,nT,nA,nG,nT,nG,nC,nG,nA,nG};
            len1 = 12'd1024;
            len2 = 13'd1536;

            // seq1 = '{M, A,T,G,T,P,T,F,T,Q,T,A,T,F,E,A,H,I,S,G,P,L,Q,S,V,V,V,L,E,G,S,F,P,V,P,E,V,S,W,F,R,D,G,Q,V,I,S,T,S,T,L,P,G,V,Q,I,S,F,S,D,G,R,A,K,L,T,I,P,A,V,T,K,A,N,S,G,R,Y,S,L,K,A,T,N,G,S,G,Q,A,T,S,T,A,E,L,L,V,K,A,E,T,A,P,P,N,F,V,Q,R,L,Q,S,M,T,V,R,Q,G,S,Q,V,R,L,Q,V,R,V,T,G,I,P,T,P,V,V,K,F,Y,R,D,G,A,E,I,Q,S,S,L,D,F,Q,I,S,Q,E,G,D,L,Y,S,L,L,I,A,E,A,Y,P,E,D,S,G,T,Y,S,V,N,A,T,N,S,V,G,R,A,T,S,T,A,E,L,L,V,Q,G,E,E,E,V,P,A,K,K,T,K,T,I,V,S,T,A,Q,I,S,E,S,R,Q,T,R,I,E,K,K,I,E,A,H,F,D,A,R,S,I,A,T,V,E,M,V,I,D,G,A,A,G,Q,Q,L,P,H,K,T,P,P,R,I,P,P,K,P,K,S,R,S,P,T,P,P,S,I,A,A,K,A,Q,L,A,R,Q,Q,S,P,S,P,I,R,H,S,P,S,P,V,R,H,V,R,A,P,T,P,S,P,V,R,S,V,S,P,A,A,R,I,S,T,S,P,I,R,S,V,R,S,P,L,L,M,R,K,T,Q,A,S,T,V,A,T,G,P,E,V,P,P,P,W,K,Q,E,G,Y,V,A,S,S,S,E,A,E,M,R,E,T,T,L,T,T,S,T,Q,I,R,T,E,E,R,W,E,G,R,Y,G,V,Q,E,Q,V,T,I,S,G,A,A,G,A,A,A,S,V,S,A,S,A,S,Y,A,A,E,A,V,A,T,G,A,K,E,V,K,Q,D,A,D,K,S,A,A,V,A,T,V,V,A,A,V,D,M,A,R,V,R,E,P,V,I,S,A,V,E,Q,T,A,Q,R,T,T,T,T,A,V,H,I,Q,P,A,Q,E,Q,V,R,K,E,A,E,K,T,A,V,T,K,V,V,V,A,A,D,K,A,K,E,Q,E,L,K,S,R,T,K,E,V,I,T,T,K,Q,E,Q,M,H,V,T,H,E,Q,I,R,K,E,T,E,K,T,F,V,P,K,V,V,I,S,A,A,K,A,K,E,Q,E,T,R,I,S,E,E,I,T,K,K,Q,K,Q,V,T,Q,E,A,I,R,Q,E,T,E,I,T,A,A,S,M,V,V,V,A,T,A,K,S,T,K,L,E,T,V,P,G,A,Q,E,E,T,T,T,Q,Q,D,Q,M,H,L,S,Y,E,K,I,M,K,E,T,R,K,T,V,V,P,K,V,I,V,A,T,P,K,V,K,E,Q,D,L,V,S,R,G,R,E,G,I,T,T,K,R,E,Q,V,Q,I,T,Q,E,K,M,R,K,E,A,E,K,T,A,L,S,T,I,A,V,A,T,A,K,A,K,E,Q,E,T,I,L,R,T,R,E,T,M,A,T,R,Q,E,Q,I,Q,V,T,H,G,K,V,D,V,G,K,K,A,E,A,V,A,T,V,V,A,A,V,D,Q,A,R,V,R,E,P,R,E,P,G,H,L,E,E,S,Y,A,Q,Q,T,T,L,E,Y,G,Y,K,E,R,I,S,A,A,K,V,A,E,P,P,Q,R,P,A,S,E,P,H,V,V,P,K,A,V,K,P,R,V,I,Q,A,P,S,E,T,H,I,K,T,T,D,Q,K,G,M,H,I,S,S,Q,I,K,K,T,T,D,L,T,T,E,R,L,V,H,V,D,K,R,P,R,T,A,S,P,H,F,T,V,S,K,I,S,V,P,K,T,E,H,G,Y,E,A,S,I,A,G,S,A,I,A,T,L,Q,K,E,L,S,A,T,S,S,A,Q,K,I,T,K,S,V,K,A,P,T,V,K,P,S,E,T,R,V,R,A,E,P,T,P,L,P,Q,F,P,F,A,D,T,P,D,T,Y,K,S,E,A,G,V,E,V,K,K,E,V,G,V,S,I,T,G,T,T,V,R,E,E,R,F,E,V,L,H,G,R,E,A,K,V,T,E,T,A,R,V,P,A,P,V,E,I,P,V,T,P,P,T,L,V,S,G,L,K,N,V,T,V,I,E,G,E,S,V,T,L,E,C,H,I,S,G,Y,P,S,P,T,V,T,W,Y,R,E,D,Y,Q,I,E,S,S,I,D,F,Q,I,T,F,Q,S,G,I,A,R,L,M,I,R,E,A,F,A,E,D,S,G,R,F,T,C,S,A,V,N,E,A,G,T,V};
            // seq2 = '{M, T,A,G,T,L,Q,S,V,V,V,L,E,G,S,T,A,T,P,M,F,T,Q,P,F,E,A,H,V,S,G,S,P,V,P,E,V,S,W,F,R,D,G,Q,V,I,S,T,S,T,L,P,G,V,Q,I,S,F,S,D,G,R,A,R,L,M,I,P,A,V,T,K,A,N,S,G,R,Y,S,L,R,A,T,N,G,S,G,Q,A,T,S,T,A,E,L,L,V,T,A,E,T,A,P,P,N,F,S,Q,R,L,Q,S,M,T,V,R,Q,G,S,Q,V,R,L,Q,V,R,V,T,G,I,P,T,P,V,V,K,F,Y,R,D,G,A,E,I,Q,S,S,L,D,F,Q,I,S,Q,E,G,D,L,Y,S,L,L,I,A,E,A,Y,P,E,D,S,G,T,Y,S,V,N,A,T,N,S,V,G,R,A,T,S,T,A,E,L,V,V,Q,G,E,E,V,V,P,A,K,K,T,K,T,I,V,S,T,A,Q,I,S,E,T,R,Q,T,R,I,E,K,K,I,E,A,H,F,D,A,R,S,I,A,T,V,E,M,V,I,D,G,A,T,G,Q,L,P,H,K,T,P,P,R,I,P,P,K,P,K,S,R,S,P,T,P,P,S,I,A,A,K,A,Q,L,A,R,Q,Q,S,P,S,P,I,R,H,S,P,S,P,V,R,H,V,R,A,P,T,P,S,P,V,R,S,V,S,P,A,G,R,I,S,T,S,P,I,R,S,V,K,S,P,L,L,I,R,K,T,Q,T,T,T,M,A,T,G,P,E,V,P,P,P,W,K,Q,E,G,Y,V,A,S,S,T,E,A,E,M,R,E,T,T,M,T,S,S,T,Q,I,R,R,E,E,R,W,E,G,R,Y,G,V,Q,E,Q,V,T,I,S,G,A,A,A,A,A,A,S,A,S,V,S,S,S,F,T,A,G,A,I,T,T,G,T,K,E,V,K,Q,E,T,D,K,S,A,A,V,A,T,V,V,A,A,V,D,M,A,R,V,R,E,P,A,I,S,A,V,E,Q,T,A,Q,R,T,T,T,T,A,V,H,I,Q,P,A,Q,E,Q,A,R,K,E,A,E,K,T,A,V,T,K,V,V,V,A,A,D,K,A,K,E,Q,E,L,K,S,R,T,R,E,V,M,V,T,T,Q,E,Q,T,H,I,S,H,E,Q,I,R,K,E,T,E,K,A,F,V,P,K,V,V,I,S,A,T,K,A,K,E,Q,E,T,R,I,T,G,E,I,T,T,K,Q,E,Q,K,R,I,T,Q,E,T,I,R,Q,E,T,E,E,I,A,A,S,M,V,V,V,A,T,A,K,S,T,K,L,E,A,A,V,G,V,Q,E,E,T,A,I,Q,Q,D,Q,M,H,L,T,H,E,Q,M,M,K,E,T,R,K,T,V,V,P,K,V,I,V,A,T,P,K,I,K,E,Q,D,L,V,S,R,S,R,E,A,I,T,T,K,R,D,Q,V,Q,I,T,Q,E,K,K,R,K,E,V,E,T,T,A,L,S,T,I,A,V,A,T,A,K,A,K,E,Q,E,T,V,L,R,S,R,E,A,M,A,T,R,Q,E,H,I,Q,V,T,H,G,Q,V,G,V,G,K,K,A,E,A,V,A,T,V,V,A,A,V,D,Q,A,R,V,R,E,P,R,E,P,T,H,V,E,E,S,H,S,Q,Q,T,T,L,E,Y,G,Y,K,E,H,I,S,T,T,K,V,P,E,Q,P,R,R,P,A,S,E,P,H,V,V,P,Q,A,V,K,P,A,V,I,Q,A,P,S,E,T,H,I,K,T,T,D,Q,M,G,M,H,I,S,S,Q,V,K,K,T,T,D,I,S,T,E,R,L,V,H,V,D,K,R,P,R,T,A,S,P,H,F,T,V,S,K,I,S,V,P,K,T,E,H,G,Y,E,A,S,I,A,G,S,A,I,A,T,L,Q,K,E,L,S,A,T,S,S,T,Q,K,I,T,K,S,V,K,A,P,T,V,K,P,G,E,T,R,V,R,A,E,P,T,P,S,P,Q,F,P,F,A,D,M,P,P,P,D,T,Y,K,S,Q,A,G,I,E,V,K,K,E,V,G,V,S,I,S,G,S,T,V,R,E,E,H,F,E,V,L,R,G,R,E,A,K,V,T,E,T,A,R,V,P,A,P,A,E,V,P,V,T,P,P,T,L,V,S,G,L,K,N,V,T,V,I,E,G,E,S,V,T,L,E,C,H,I,S,G,Y,P,S,P,K,V,T,W,Y,R,E,D,Y,Q,I,E,S,S,I,D,F,Q,I,T,F,Q,G,G,I,A,R,L,M,I,R,E,A,F,A,E,D,S,G,R,F,T,C,S,A,V,N,E,A};
            // len1 = 12'd5;
            // len2 = 12'd5;
            // seq1 = '{M, T,T,Q,A,P,T,F,T,Q,T,A,T,F,E,A,H,I,S,G,P,L,Q,S,V,V,V,L,E,G,S,F,P,V,P,E,V,S,W,F,R,D,G,Q,V,I,S,T,S,T,L,P,G,V,Q,I,S,F,S,D,G,R,A,K,L,T,I,P,A,V,T,K,A,N,S,G,R,Y,S,L,K,A,T,N,G,S,G,Q,A,T,S,T,A,E,L,L,V,K,A,E,T,A,P,P,N,F,V,Q,R,L,Q,S,M,T,V,R,Q,G,S,Q,V,R,L,Q,V,R,V,T,G,I,P,T,P,V,V,K,F,Y,R,D,G,A,E,I,Q,S,S,L,D,F,Q,I,S,Q,E,G,D,L,Y,S,L,L,I,A,E,A,Y,P,E,D,S,G,T,Y,S,V,N,A,T,N,S,V,G,R,A,T,S,T,A,E,L,L,V,Q,G,E,E,E,V,P,A,K,K,T,K,T,I,V,S,T,A,Q,I,S,E,S,R,Q,T,R,I,E,K,K,I,E,A,H,F,D,A,R,S,I,A,T,V,E,M,V,I,D,G,A,A,G,Q,Q,L,P,H,K,T,P,P,R,I,P,P,K,P,K,S,R,S,P,T,P,P,S,I,A,A,K,A,Q,L,A,R,Q,Q,S,P,S,P,I,R,H,S,P,S,P,V,R,H,V,R,A,P,T,P,S,P,V,R,S,V,S,P,A,A,R,I,S,T,S,P,I,R,S,V,R,S,P,L,L,M,R,K,T,Q,A,S,T,V,A,T,G,P,E,V,P,P,P,W,K,Q,E,G,Y,V,A,S,S,S,E,A,E,M,R,E,T,T,L,T,T,S,T,Q,I,R,T,E,E,R,W,E,G,R,Y,G,V,Q,E,Q,V,T,I,S,G,A,A,G,A,A,A,S,V,S,A,S,A,S,Y,A,A,E,A,V,A,T,G,A,K,E,V,K,Q,D,A,D,K,S,A,A,V,A,T,V,V,A,A,V,D,M,A,R,V,R,E,P,V,I,S,A,V,E,Q,T,A,Q,R,T,T,T,T,A,V,H,I,Q,P,A,Q,E,Q,V,R,K,E,A,E,K,T,A,V,T,K,V,V,V,A,A,D,K,A,K,E,Q,E,L,K,S,R,T,K,E,V,I,T,T,K,Q,E,Q,M,H,V,T,H,E,Q,I,R,K,E,T,E,K,T,F,V,P,K,V,V,I,S,A,A,K,A,K,E,Q,E,T,R,I,S,E,E,I,T,K,K,Q,K,Q,V,T,Q,E,A,I,R,Q,E,T,E,I,T,A,A,S,M,V,V,V,A,T,A,K,S,T,K,L,E,T,V,P,G,A,Q,E,E,T,T,T,Q,Q,D,Q,M,H,L,S,Y,E,K,I,M,K,E,T,R,K,T,V,V,P,K,V,I,V,A,T,P,K,V,K,E,Q,D,L,V,S,R,G,R,E,G,I,T,T,K,R,E,Q,V,Q,I,T,Q,E,K,M,R,K,E,A,E,K,T,A,L,S,T,I,A,V,A,T,A,K,A,K,E,Q,E,T,I,L,R,T,R,E,T,M,A,T,R,Q,E,Q,I,Q,V,T,H,G,K,V,D,V,G,K,K,A,E,A,V,A,T,V,V,A,A,V,D,Q,A,R,V,R,E,P,R,E,P,G,H,L,E,E,S,Y,A,Q,Q,T,T,L,E,Y,G,Y,K,E,R,I,S,A,A,K,V,A,E,P,P,Q,R,P,A,S,E,P,H,V,V,P,K,A,V,K,P,R,V,I,Q,A,P,S,E,T,H,I,K,T,T,D,Q,K,G,M,H,I,S,S,Q,I,K,K,T,T,D,L,T,T,E,R,L,V,H,V,D,K,R,P,R,T,A,S,P,H,F,T,V,S,K,I,S,V,P,K,T,E,H,G,Y,E,A,S,I,A,G,S,A,I,A,T,L,Q,K,E,L,S,A,T,S,S,A,Q,K,I,T,K,S,V,K,A,P,T,V,K,P,S,E,T,R,V,R,A,E,P,T,P,L,P,Q,F,P,F,A,D,T,P,D,T,Y,K,S,E,A,G,V,E,V,K,K,E,V,G,V,S,I,T,G,T,T,V,R,E,E,R,F,E,V,L,H,G,R,E,A,K,V,T,E,T,A,R,V,P,A,P,V,E,I,P,V,T,P,P,T,L,V,S,G,L,K,N,V,T,V,I,E,G,E,S,V,T,L,E,C,H,I,S,G,Y,P,S,P,T,V,T,W,Y,R,E,D,Y,Q,I,E,S,S,I,D,F,Q,I,T,F,Q,S,G,I,A,R,L,M,I,R,E,A,F,A,E,D,S,G,R,F,T,C,S,A,V,N,E,A,G,T,V};
            // seq2 = '{M, T,T,Q,A,L,Q,S,V,V,V,L,E,G,S,T,A,T,P,M,F,T,Q,P,F,E,A,H,V,S,G,S,P,V,P,E,V,S,W,F,R,D,G,Q,V,I,S,T,S,T,L,P,G,V,Q,I,S,F,S,D,G,R,A,R,L,M,I,P,A,V,T,K,A,N,S,G,R,Y,S,L,R,A,T,N,G,S,G,Q,A,T,S,T,A,E,L,L,V,T,A,E,T,A,P,P,N,F,S,Q,R,L,Q,S,M,T,V,R,Q,G,S,Q,V,R,L,Q,V,R,V,T,G,I,P,T,P,V,V,K,F,Y,R,D,G,A,E,I,Q,S,S,L,D,F,Q,I,S,Q,E,G,D,L,Y,S,L,L,I,A,E,A,Y,P,E,D,S,G,T,Y,S,V,N,A,T,N,S,V,G,R,A,T,S,T,A,E,L,V,V,Q,G,E,E,V,V,P,A,K,K,T,K,T,I,V,S,T,A,Q,I,S,E,T,R,Q,T,R,I,E,K,K,I,E,A,H,F,D,A,R,S,I,A,T,V,E,M,V,I,D,G,A,T,G,Q,L,P,H,K,T,P,P,R,I,P,P,K,P,K,S,R,S,P,T,P,P,S,I,A,A,K,A,Q,L,A,R,Q,Q,S,P,S,P,I,R,H,S,P,S,P,V,R,H,V,R,A,P,T,P,S,P,V,R,S,V,S,P,A,G,R,I,S,T,S,P,I,R,S,V,K,S,P,L,L,I,R,K,T,Q,T,T,T,M,A,T,G,P,E,V,P,P,P,W,K,Q,E,G,Y,V,A,S,S,T,E,A,E,M,R,E,T,T,M,T,S,S,T,Q,I,R,R,E,E,R,W,E,G,R,Y,G,V,Q,E,Q,V,T,I,S,G,A,A,A,A,A,A,S,A,S,V,S,S,S,F,T,A,G,A,I,T,T,G,T,K,E,V,K,Q,E,T,D,K,S,A,A,V,A,T,V,V,A,A,V,D,M,A,R,V,R,E,P,A,I,S,A,V,E,Q,T,A,Q,R,T,T,T,T,A,V,H,I,Q,P,A,Q,E,Q,A,R,K,E,A,E,K,T,A,V,T,K,V,V,V,A,A,D,K,A,K,E,Q,E,L,K,S,R,T,R,E,V,M,V,T,T,Q,E,Q,T,H,I,S,H,E,Q,I,R,K,E,T,E,K,A,F,V,P,K,V,V,I,S,A,T,K,A,K,E,Q,E,T,R,I,T,G,E,I,T,T,K,Q,E,Q,K,R,I,T,Q,E,T,I,R,Q,E,T,E,E,I,A,A,S,M,V,V,V,A,T,A,K,S,T,K,L,E,A,A,V,G,V,Q,E,E,T,A,I,Q,Q,D,Q,M,H,L,T,H,E,Q,M,M,K,E,T,R,K,T,V,V,P,K,V,I,V,A,T,P,K,I,K,E,Q,D,L,V,S,R,S,R,E,A,I,T,T,K,R,D,Q,V,Q,I,T,Q,E,K,K,R,K,E,V,E,T,T,A,L,S,T,I,A,V,A,T,A,K,A,K,E,Q,E,T,V,L,R,S,R,E,A,M,A,T,R,Q,E,H,I,Q,V,T,H,G,Q,V,G,V,G,K,K,A,E,A,V,A,T,V,V,A,A,V,D,Q,A,R,V,R,E,P,R,E,P,T,H,V,E,E,S,H,S,Q,Q,T,T,L,E,Y,G,Y,K,E,H,I,S,T,T,K,V,P,E,Q,P,R,R,P,A,S,E,P,H,V,V,P,Q,A,V,K,P,A,V,I,Q,A,P,S,E,T,H,I,K,T,T,D,Q,M,G,M,H,I,S,S,Q,V,K,K,T,T,D,I,S,T,E,R,L,V,H,V,D,K,R,P,R,T,A,S,P,H,F,T,V,S,K,I,S,V,P,K,T,E,H,G,Y,E,A,S,I,A,G,S,A,I,A,T,L,Q,K,E,L,S,A,T,S,S,T,Q,K,I,T,K,S,V,K,A,P,T,V,K,P,G,E,T,R,V,R,A,E,P,T,P,S,P,Q,F,P,F,A,D,M,P,P,P,D,T,Y,K,S,Q,A,G,I,E,V,K,K,E,V,G,V,S,I,S,G,S,T,V,R,E,E,H,F,E,V,L,R,G,R,E,A,K,V,T,E,T,A,R,V,P,A,P,A,E,V,P,V,T,P,P,T,L,V,S,G,L,K,N,V,T,V,I,E,G,E,S,V,T,L,E,C,H,I,S,G,Y,P,S,P,K,V,T,W,Y,R,E,D,Y,Q,I,E,S,S,I,D,F,Q,I,T,F,Q,G,G,I,A,R,L,M,I,R,E,A,F,A,E,D,S,G,R,F,T,C,S,A,V,N,E,A};
            // len1 = 12'd53;
            // len2 = 12'd53;

            #20 rst = 0; // after 2 clock ticks set reset to inactive (0)

            #5 wrreq = 1'b1;
            wren = 1'b1;
            #10 in16 = 16'hF0F0;
            wraddress = 15'd3;
            in2 = 2'b01;

            solver_enable = 1;

            #10 wrreq = 1'b0;
            wren = 1'b0;
            #10 rdreq = 1'b1;
            rdaddress = 15'd3;

            #40 rdreq = 1'b0;

            // #12000 rst = 1;
            // solver_enable = 0;

            // seq1 = '{nA, nA,nG,nG,nA,nG,nG,nG,nG,nG,nC,nG,nT,nT,nG,nA,nT,nG,nT,nG,nG,nC,nC,nG,nT,nC,nT,nG,nT,nT,nT,nG,nT,nG,nA,nC,nG,nT,nA,nT,nG,nT,nA,nG,nA,nC,nA,nG,nC,nA,nA,nC,nG,nC,nT,nC,nT,nC,nT,nC,nA,nG,nC,nC,nC,nT,nG,nT,nT,nG,nT,nT,nG,nT,nC,nT,nC,nT,nA,nT,nC,nC,nA,nA,nC,nC,nC,nC,nG,nG,nC,nC,nC,nT,nA,nT,nA,nA,nA,nT,nT,nT,nT,nT,nG,nA,nG,nA,nT,nG,nT,nC,nC,nG,nA,nC,nG,nA,nC,nC,nG,nG,nT,nC,nA,nG,nA,nA,nA,nT,nC,nC,nT,nG,nG,nT,nT,nC,nA,nG,nC,nG,nC,nA,nA,nA,nA,nG,nG,nT,nC,nA,nC,nT,nT,nA,nA,nG,nA,nT,nC,nA,nA,nA,nG,nA,nA,nG,nG,nG,nG,nC,nA,nC,nC,nA,nT,nC,nC,nG,nA,nG,nT,nT,nT,nC,nC,nC,nT,nT,nC,nT,nG,nA,nA,nG,nT,nA,nG,nT,nT,nC,nT,nT,nC,nC,nA,nG,nA,nT,nC,nT,nT,nC,nT,nT,nG,nC,nT,nC,nC,nG,nA,nC,nA,nT,nA,nC,nA,nG,nT,nC,nG,nA,nA,nG,nG,nG,nA,nT,nA,nA,nT,nA,nC,nC,nA,nT,nC,nA,nA,nC,nT,nA,nG,nC,nG,nT,nC,nA,nA,nC,nT,nC,nA,nA,nC,nT,nC,nA,nC,nT,nG,nG,nT,nA,nG,nT,nT,nC,nC,nT,nG,nC,nT,nG,nA,nG,nA,nA,nT,nA,nC,nT,nT,nT,nA,nT,nA,nT,nG,nT,nG,nA,nA,nA,nT,nG,nG,nC,nA,nT,nG,nC,nC,nA,nT,nA,nG,nT,nA,nC,nT,nG,nC,nA,nC,nC,nA,nA,nG,nC,nG,nC,nT,nG,nA,nA,nT,nT,nA,nG,nT,nA,nT,nC,nG,nG,nA,nT,nG,nG,nT,nA,nT,nT,nC,nA,nG,nC,nA,nT,nG,nC,nC,nT,nA,nA,nA,nG,nG,nC,nA,nT,nG,nG,nG,nT,nT,nA,nC,nC,nT,nC,nG,nC,nC,nC,nG,nG,nT,nT,nA,nC,nC,nT,nA,nC,nG,nC,nA,nT,nT,nA,nG,nA,nC,nT,nG,nG,nT,nC,nA,nT,nA,nG,nA,nC,nC,nC,nC,nG,nT,nA,nT,nT,nA,nT,nC,nT,nT,nT,nT,nC,nT,nC,nT,nG,nG,nG,nC,nC,nA,nC,nG,nC,nA,nG,nG,nC,nT,nG,nT,nT,nC,nA,nC,nC,nG,nC,nT,nG,nA,nG,nC,nG,nG,nT,nC,nG,nA,nC,nA,nC,nC,nG,nA,nT,nG,nC,nT,nG,nG,nA,nG,nG,nG,nT,nT,nG,nC,nG,nA,nG,nC,nA,nC,nG,nT,nA,nG,nC,nA,nG,nG,nC,nA,nT,nC,nA,nT,nC,nT,nG,nG,nA,nC,nA,nG,nT,nG,nG,nG,nT,nA,nA,nG,nA,nT,nT,nA,nC,nG,nG,nC,nT,nT,nA,nA,nT,nT,nG,nT,nA,nT,nC,nG,nC,nG,nT,nC,nG,nG,nA,nA,nC,nG,nA,nA,nC,nA,nA,nG,nG,nT,nG,nC,nA,nG,nC,nA,nT,nA,nT,nC,nC,nG,nT,nA,nA,nT,nT,nT,nT,nC,nT,nC,nC,nA,nA,nA,nT,nC,nG,nC,nA,nC,nC,nA,nT,nT,nG,nG,nA,nA,nC,nA,nG,nC,nT,nA,nA,nA,nG,nT,nG,nA,nG,nA,nG,nA,nA,nC,nC,nG,nT,nA,nG,nG,nT,nA,nT,nC,nC,nC,nT,nC,nA,nC,nG,nG,nA,nC,nC,nG,nC,nC,nA,nC,nC,nA,nA,nA,nT,nC,nA,nA,nA,nA,nC,nC,nT,nT,nA,nA,nA,nC,nG,nT,nA,nT,nG,nG,nC,nA,nT,nT,nA,nG,nG,nC,nT,nA,nA,nC,nC,nA,nC,nA,nC,nT,nT,nA,nG,nT,nC,nA,nT,nG,nG,nC,nC,nG,nC,nG,nT,nT,nC,nC,nT,nG,nG,nA,nC,nG,nA,nG,nG,nG,nA,nC,nG,nG,nA,nA,nA,nT,nT,nA,nA,nG,nG,nG,nC,nC,nG,nT,nG,nG,nA,nG,nG,nG,nA,nC,nC,nC,nT,nG,nG,nC,nG,nA,nC,nA,nG,nG,nT,nC,nT,nA,nA,nC,nG,nG,nG,nT,nG,nT,nT,nC,nC,nT,nA,nT,nA,nT,nC,nC,nA,nA,nC,nC,nT,nC,nT,nA,nG,nC,nA,nT,nC,nC,nC,nT,nA,nC,nA,nC,nG,nT,nA,nG,nA,nC,nC,nT,nC,nA,nA,nT,nG,nA,nG,nC,nG,nG,nT,nG,nC,nG,nC,nA,nA,nG,nA,nT,nT,nT,nG,nC,nC,nC,nT,nT,nA,nG,nA,nT,nG,nT,nG,nC,nG,nC,nT,nC,nA,nT,nG,nC,nT,nT,nT,nG,nT,nC,nT,nT,nT,nA,nG,nA,nC,nC,nC,nC,nG,nA,nA,nC,nT,nC,nT,nG,nC,nA,nG,nG,nC,nT,nC,nC,nA,nC,nA,nT,nC,nT,nG,nT,nT,nT,nC,nA,nC,nG,nA,nT,nA,nA,nA,nT,nC,nC,nC,nA,nG,nC,nG,nT,nC,nT,nA,nT,nG,nA,nT,nG,nT,nG,nG,nT,nA,nG,nC,nG,nT,nC,nC,nC,nG,nT,nC,nA,nT,nC,nT,nA,nT,nT,nA,nC,nG,nG,nT,nA,nA,nT,nG,nG,nC,nC,nG,nT,nT,nA,nT,nG,nA,nA,nT,nG,nT,nC,nT,nT,nA,nT,nG,nC,nT,nG,nC,nC,nG,nA,nG,nC,nT,nT,nC,nT,nG,nG,nA,nC,nG,nA,nG,nT,nC,nT,nA,nG,nT,nC,nT,nC,nC,nT,nA,nT,nA,nG,nT,nA,nT,nG,nG,nG,nA,nC,nG,nG,nG,nC,nT,nC,nT,nG,nA,nC,nT};
            // seq2 = '{nA, nG,nG,nC,nT,nG,nC,nG,nT,nC,nT,nT,nC,nA,nA,nC,nG,nA,nC,nC,nT,nT,nT,nC,nA,nC,nC,nT,nT,nT,nG,nC,nA,nT,nC,nT,nC,nG,nA,nC,nG,nA,nA,nT,nT,nT,nC,nG,nA,nT,nC,nG,nT,nA,nT,nG,nG,nA,nT,nA,nT,nT,nC,nT,nA,nC,nC,nG,nA,nG,nT,nT,nG,nC,nC,nA,nT,nG,nG,nA,nC,nG,nG,nG,nG,nA,nA,nC,nG,nA,nG,nT,nG,nG,nA,nT,nA,nC,nA,nC,nC,nT,nC,nC,nC,nG,nA,nC,nT,nT,nT,nA,nA,nA,nC,nA,nG,nA,nA,nA,nT,nC,nG,nT,nC,nG,nC,nA,nT,nA,nC,nT,nC,nT,nG,nC,nC,nT,nA,nT,nC,nG,nC,nA,nC,nT,nC,nT,nT,nG,nA,nC,nT,nA,nC,nA,nT,nG,nG,nT,nG,nG,nG,nG,nA,nC,nT,nC,nC,nT,nT,nA,nT,nC,nA,nG,nC,nT,nC,nG,nA,nC,nT,nT,nG,nG,nG,nG,nC,nC,nC,nA,nA,nG,nG,nT,nA,nC,nA,nA,nG,nT,nA,nG,nG,nT,nT,nG,nA,nA,nA,nC,nG,nG,nC,nC,nC,nG,nG,nC,nG,nT,nT,nG,nT,nT,nG,nG,nC,nG,nT,nC,nA,nC,nT,nC,nT,nT,nA,nG,nC,nA,nC,nA,nC,nT,nG,nA,nC,nG,nC,nT,nC,nC,nT,nA,nG,nC,nT,nG,nA,nG,nA,nC,nC,nT,nT,nG,nA,nA,nC,nA,nT,nG,nC,nA,nG,nG,nA,nC,nG,nT,nC,nC,nC,nT,nG,nT,nG,nC,nC,nA,nA,nT,nT,nC,nG,nC,nT,nA,nT,nG,nG,nG,nC,nC,nT,nT,nC,nA,nA,nG,nG,nA,nT,nT,nT,nC,nA,nT,nA,nG,nC,nA,nT,nT,nA,nC,nC,nG,nT,nC,nT,nC,nA,nC,nG,nG,nC,nC,nA,nC,nG,nC,nA,nG,nG,nG,nC,nG,nC,nG,nA,nT,nG,nA,nA,nC,nC,nC,nG,nG,nT,nT,nA,nG,nT,nT,nG,nA,nT,nT,nT,nT,nG,nT,nG,nA,nT,nT,nT,nA,nT,nT,nT,nC,nG,nT,nG,nT,nG,nG,nT,nC,nA,nT,nA,nC,nG,nC,nG,nG,nA,nT,nT,nC,nT,nT,nA,nC,nT,nA,nA,nG,nT,nC,nT,nC,nT,nA,nC,nG,nG,nA,nA,nG,nA,nA,nC,nC,nC,nT,nC,nG,nA,nT,nA,nG,nG,nA,nG,nT,nC,nC,nG,nA,nC,nA,nA,nT,nG,nG,nA,nG,nA,nA,nT,nA,nA,nC,nT,nA,nA,nA,nG,nA,nA,nG,nC,nG,nC,nT,nT,nC,nG,nA,nC,nC,nC,nC,nA,nA,nG,nC,nG,nA,nC,nA,nG,nC,nG,nA,nA,nT,nC,nG,nG,nG,nA,nT,nT,nT,nG,nC,nG,nA,nG,nA,nA,nC,nT,nC,nA,nC,nA,nG,nG,nA,nT,nC,nC,nA,nT,nC,nA,nA,nG,nT,nC,nC,nT,nA,nC,nC,nG,nT,nC,nG,nC,nT,nG,nA,nG,nC,nA,nG,nG,nT,nC,nC,nT,nG,nG,nG,nA,nC,nA,nG,nT,nA,nG,nT,nT,nC,nC,nA,nG,nT,nT,nA,nT,nT,nC,nC,nT,nA,nA,nT,nA,nG,nA,nC,nT,nC,nA,nG,nC,nT,nC,nC,nA,nG,nC,nA,nG,nG,nA,nG,nC,nG,nA,nC,nT,nA,nA,nA,nA,nG,nG,nT,nC,nA,nA,nA,nG,nG,nG,nA,nC,nC,nT,nC,nT,nT,nG,nG,nG,nG,nT,nT,nG,nA,nG,nC,nG,nA,nC,nC,nT,nG,nT,nG,nT,nT,nT,nT,nA,nA,nC,nG,nC,nC,nA,nG,nG,nC,nC,nC,nT,nA,nA,nC,nC,nC,nC,nG,nC,nC,nT,nG,nG,nA,nG,nG,nG,nC,nC,nC,nG,nC,nA,nA,nG,nT,nG,nG,nT,nC,nA,nG,nC,nT,nG,nT,nT,nC,nT,nA,nG,nT,nA,nC,nA,nG,nT,nT,nA,nC,nT,nG,nA,nT,nC,nA,nG,nA,nA,nT,nC,nA,nC,nT,nG,nT,nC,nC,nG,nC,nC,nT,nA,nC,nC,nC,nG,nT,nT,nC,nA,nT,nC,nC,nA,nA,nC,nG,nT,nG,nG,nT,nT,nT,nG,nA,nC,nG,nA,nT,nT,nC,nC,nC,nG,nA,nG,nG,nG,nT,nA,nA,nT,nA,nT,nA,nG,nG,nC,nC,nG,nG,nC,nA,nC,nT,nA,nT,nT,nC,nG,nC,nG,nG,nC,nG,nT,nT,nA,nG,nT,nT,nG,nT,nT,nC,nT,nT,nC,nC,nT,nG,nC,nC,nG,nG,nA,nC,nA,nC,nC,nT,nA,nT,nC,nC,nT,nC,nG,nA,nC,nT,nC,nG,nG,nC,nG,nC,nG,nG,nG,nG,nA,nG,nC,nC,nA,nG,nA,nA,nC,nG,nC,nG,nA,nT,nG,nT,nG,nT,nG,nA,nA,nC,nT,nT,nC,nG,nG,nT,nC,nC,nG,nG,nC,nA,nA,nA,nA,nA,nA,nA,nC,nC,nA,nT,nA,nT,nC,nG,nT,nG,nG,nT,nA,nC,nC,nG,nC,nT,nA,nG,nT,nA,nA,nT,nC,nA,nC,nT,nT,nC,nT,nA,nG,nT,nT,nT,nC,nT,nG,nT,nG,nA,nA,nG,nT,nC,nG,nG,nA,nC,nT,nC,nC,nG,nA,nT,nC,nC,nG,nA,nA,nC,nC,nA,nA,nG,nA,nG,nT,nA,nC,nG,nG,nA,nG,nA,nA,nT,nT,nC,nG,nA,nA,nG,nC,nG,nC,nT,nG,nC,nC,nG,nA,nT,nG,nC,nA,nC,nT,nC,nG,nC,nC,nA,nG,nA,nG,nG,nT,nA,nG,nC,nC,nG,nC,nA,nC,nT,nA,nA,nT,nA,nT,nC,nC,nG,nG,nT,nG,nA,nA,nC,nA,nG,nG,nT,nA,nG,nT,nG,nC,nG,nA,nG};
            // len1 = 12'd53;
            // len2 = 12'd53;

            // #20 rst = 0;
            // #10 solver_enable = 1;


        end

    always #5       // every five simulation units...
        clk <= !clk;  // ...invert the clock

                    // produce debug output on the negative edge of the clock

endmodule // tb_short_solver
